
module mvm_noc_top (
	clk_clk,
	leds_leds);	

	input		clk_clk;
	output	[9:0]	leds_leds;
endmodule
